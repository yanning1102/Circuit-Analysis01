
vcc 1 0 dc 15v
rb1 1 2 100k
rb2 2 0 50k
rc 1 3 4k
re 4 0 3k
q1 3 2 4 aaa
.model aaa npn(level=1 bf=100 is=1.8e-15a )
.op
.probe
.end