
vi 1 0 sin(0v 5v 100hz)
vb 3 0 dc -5v
vg 2 0 dc 5v
rl 4 0 100k
m1 1 2 4 3 aaa l=10u w=50u
.model aaa nmos(kp=20u vto=1v lambda=0)
.tran 0.01ms 40ms 0ms 0.01ms
.probe
.end