
vi 1 0 dc 2.4v
vbn 3 0 dc -5v
vgn 2 0 dc 5v
m1 1 2 0 3 aaa (l=10u w=50u)
.model aaa nmos(kp=20u vto=1v lambd=0)

vbp 4 0 dc 5v
vgp 5 0 dc -5v
m2 1 5 0 4 ccc(l=10u w=50u)
.model ccc pmos(kp=20u vto=1v lambd=0)
.dc vi -5 5 0.01
.probe
.end