
vdd 1 0 dc 12v
ro 1 4 200000
m3 1 1 2 0 aaa3 
m2 2 2 3 0 aaa2
m1 3 3 0 0 aaa1
m4 4 3 0 0 aaa4
.model aaa1 nmos(kp=1.073u vto=1.73 phi=0.6 gamma=0.5 lambda=0 l=240u w=2000u)
.model aaa2 nmos(kp=1.073u vto=1.73 phi=0.6 gamma=0.5 lambda=0 l=12u w=2000u)
.model aaa3 nmos(kp=1.073u vto=1.73 phi=0.6 gamma=0.5 lambda=0 l=32u w=2000u)
.model aaa4 nmos(kp=1.073u vto=1.73 phi=0.6 gamma=0.5 lambda=0 l=240u w=2000u)


.op
.probe
.end