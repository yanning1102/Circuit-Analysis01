* circuit description *
Vcc 1 0 DC 15
Vo 3 0 DC 5
RE 4 0 5k
is 1 2 dc 0.73m
*BJT model description
Q1 2 2 0 0 npn_transistor
Q2 3 2 4 0 npn_transistor

.model npn_transistor npn (Is=1.8E-15 BF=100 VAF=100)
*analysis requests
.DC Vo 0 15 0.01
*output requests
.op
.plot DC I(Vo)
.probe
.end