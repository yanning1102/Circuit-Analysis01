
*r1 1 2 11.81272234k
i1 1 2 dc 1m
vdd 1 0 dc 15
vo 3 0 dc 7
M1 2 4 0 0 e_mos L=10u W=100u
M2 4 4 0 0 e_mos L=10u W=100u
*M3 2 2 3 0 e_mos L=5u W=50u
M4 3 2 4 4 e_mos L=10u W=100u
.model e_mos nmos (KP=20u Vto=1V lambda=0.02)

.dc vo 0 15 0.1
.op
.probe
.end
