
vdd vdd 0 dc 12
*vi vi 0 sin(0 0.05 100)
vi vi 0 dc 6
M1 1 1 0 0 e_mos L=1u W=1.6322548u
M2 2 2 1 0 e_mos L=1u W=18.4516948u
M3 vdd vdd 2 0 e_mos L=1u W=18.4516948u
*M4 3 1 0 0 e_mos L=1u W=1.01u
*M5 3 vi vdd vdd d_mos L=1u W=0.31057841u
M4 3 1 0 0 e_mos L=1u W=1.01016892u
M5 3 vi vdd vdd d_mos L=1u W=0.31057841u

.model e_mos nmos (KP=1.073u Vto=1.73 lambda=0.002)
.model d_mos pmos (KP=10.43u Vto=-3.533 lambda=0.002)
.op
*.tran 0.1m 40m 0m 0.01m
.probe
.end
