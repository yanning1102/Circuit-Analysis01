
v1 2 0 dc 5
v2 3 0 dc -5
v3 4 0 dc 5
v4 5 0 dc -5

vi 1 0 dc 0

M1 1 2 0 3 e_mos L=5u W=50u
M2 1 5 0 4 s_mos L=5u W=50u

.model e_mos nmos (KP=20u Vto=2V lambda=0.02)
.model s_mos pmos (KP=20u Vto=2V lambda=0.02)
.dc vi -5 5 0.01
.op

.probe
.end
