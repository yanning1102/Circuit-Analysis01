
vdd vdd 0 dc 12
*v1 v1 0 dc 3
*v2 v2 0 dc 6
M1 1 1 0 0 e_mos L=1u W=0.54511354u
M2 2 2 1 0 e_mos L=1u W=1.75u
M3 vdd vdd 2 0 e_mos L=1u W=0.0732u
.model e_mos nmos (KP=1.073u Vto=1.73 gamma=0.5 lambda=0.02)

.op
.probe
.end
