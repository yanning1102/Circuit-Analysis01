
vdd 1 0 dc 12v
m3 2 2 1 1 bbb3
m2 2 2 3 0 aaa2
m1 3 3 0 0 aaa1
m4 4 2 1 1 bbb4
m5 4 2 5 0 aaa5
m6 5 6 0 0 aaa6
.model aaa1 nmos(kp=1.073u vto=1.73 gamma=0 lambda=0.02 w=6.64 l=0.1)
.model aaa2 nmos(kp=1.073u vto=1.73 phi=0.6 gamma=0.5 lambda=0.02 w=16.5 l=0.1)
.model bbb3 pmos(kp=10.43u vto=-3.533 gamma=0 lambda=0.02 w=0.69 l=0.1)
.model bbb4 pmos(kp=10.43u vto=-3.533 gamma=0 lambda=0.02 w=0.707 l=0.1)
.model aaa5 nmos(kp=1.073u vto=1.73 phi=0.6 gamma=0.5 lambda=0.02 w=5154 l=0.1)
.model aaa6 nmos(kp=1.073u vto=1.73 gamma=0 lambda=0.02 w=6.67 l=0.1)
vi 6 7 dc 3.4v
vs 7 0 sin(0 0.00334 1k 0 0 0)
.op
.tran 0.01 20m 0 0.01
.probe
.end