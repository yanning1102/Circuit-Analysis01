
vdd vdd 0 dc 12
vi vi 0 dc 3
vg vg 0 dc 6

M1 1 1 0 0 e_mos L=1u W=11.48748218u
M2 2 2 1 0 e_mos L=1u W=11.49u
M3 2 2 vdd vdd d_mos L=1u W=0.31133423u
M4 3 2 vdd vdd d_mos L=1u W=0.31133423u
M5 3 vg vi 0 e_mos L=1u W=11.4881u
.model e_mos nmos (KP=1.073u Vto=1.73 lambda=0.002)
.model d_mos pmos (KP=10.43u Vto=-3.533 lambda=0.002)
.op
.probe
.end
