

rd 3 4 4k
*rd 3 4 6k
*vdd 3 0 dc 15
vcc 3 0 dc 15
*r1 1 2 50k
*r2 2 3 20meg
*r3 3 0 20meg
vi 2 1 dc 0
vgs 1 0 dc 6
*vds 2 0 dc 0
M1 4 2 0 0 e_mos L=5u W=50u

.model e_mos nmos (KP=20u Vto=2V lambda=0.02)

.dc vi 0 15 0.01
.probe
.end
