
vcc 1 0 dc 15v
iref 1 2 dc 0.73m
q1 2 2 0 aaa
.model aaa npn(is=1.8e-15 vaf=100 bf=100)
vo 3 0 dc 5v
q2 3 2 4 bbb
.model bbb npn(is=1.8e-15 vaf=100 bf=100)
re 4 0 5k
.op
.dc vo 0 15 0.01
.plot dc i(vo)
.probe
.end