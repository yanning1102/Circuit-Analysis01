
v1 2 0 dc 5
v2 3 0 dc -5
v3 5 0 dc -5
v4 4 0 dc 5
r1 6 0 100k
*vdd 1 0 dc 10

*r1 1 2 50k
*r2 2 3 20meg
*r3 3 0 20meg
vi 1 0 sin(0 5 100 0 0 0)
M1 1 2 6 3 e_mos L=5u W=50u
M2 1 5 6 4 t_mos L=5u W=50u
.model e_mos nmos (KP=20u Vto=2V lambda=0.02)
.model t_mos pmos (KP=20u Vto=2V lambda=0.02)
.tran 0.01m 40m 0 0.01m
.probe
.end

v1 2 0 dc 5
v2 3 0 dc -5
v3 5 0 dc -5
v4 4 0 dc 5
r1 6 0 10k
*vdd 1 0 dc 10

*r1 1 2 50k
*r2 2 3 20meg
*r3 3 0 20meg
vi 1 0 sin(0 5 100 0 0 0)
M1 1 2 6 3 e_mos L=5u W=50u
M2 1 5 6 4 t_mos L=5u W=50u
.model e_mos nmos (KP=20u Vto=2V lambda=0.02)
.model t_mos pmos (KP=20u Vto=2V lambda=0.02)
.tran 0.01m 40m 0 0.01m
.probe
.end

v1 2 0 dc 5
v2 3 0 dc -5
v3 5 0 dc -5
v4 4 0 dc 5
r1 6 0 1k
*vdd 1 0 dc 10

*r1 1 2 50k
*r2 2 3 20meg
*r3 3 0 20meg
vi 1 0 sin(0 5 100 0 0 0)
M1 1 2 6 3 e_mos L=5u W=50u
M2 1 5 6 4 t_mos L=5u W=50u
.model e_mos nmos (KP=20u Vto=2V lambda=0.02)
.model t_mos pmos (KP=20u Vto=2V lambda=0.02)
.tran 0.01m 40m 0 0.01m
.probe
.end
