*circuit description
Vi 1 0 dc 0
*sin(0V 10V 60HZ)
VR1 4 0 dc 5V
VR2 6 0 dc -5V
R1 1 2 10k
R2 2 3 10k
R3 2 5 10k
*diode model descriotion
D1 3 4 1mA_diode
D2 6 5 1mA_diode
.model 1mA_diode D (Is=0.01pA n=1.0675)
*analysis requests
*.TRAN 0.01ms 40ms 0ms 0.01ms
.dc Vi -10 10 0.01
.probe
.end