
vg 2 0 dc 5
vb 3 0 dc -5
*vdd 1 0 dc 10

*r1 1 2 50k
*r2 2 3 20meg
*r3 3 0 20meg
vi 1 0 dc 0
M1 1 2 0 3 e_mos L=5u W=50u

.model e_mos nmos(KP=20u Vto=2V lambda=0.02)
.dc vi -5 5 0.01
.op

.probe
.end
