* circuit description *
Vcc 1 0 DC 15
Vo 4 0 DC 5
*R1 1 2 14.3k
is 1 2 dc 1m
*BJT model description
Q1 2 3 0 0 npn_transistor
Q2 3 3 0 0 npn_transistor
Q3 4 2 3 0 npn_transistor
.model npn_transistor npn (Is=1.8E-15 BF=100 VAF=100)
*analysis requests
.DC Vo 0 15 0.01
*output requests
.op
.plot DC I(Vo)
.probe
.end