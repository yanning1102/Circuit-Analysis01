
vi 1 0 dc 2.4v
vr1 4 0 dc 5v
vr2 6 0 dc -5v
r1 1 2 10k
r2 2 3 10k
r3 2 5 10k
d1 3 4 dio
d2 6 5 dio
.model dio d(is=0.01pa n=1.0675)
.dc vi -10 10 0.01
.probe
.end