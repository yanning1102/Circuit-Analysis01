
*circuit description
vdd vdd 0 dc 3
*vi vi 0 sin(0V 10V 60HZ)
vi vi 0 pulse(0 3 0 0 0 10u 20u)
v2 1 2 dc 0
*diode model descriotion
c1 2 0 1p
M1 1 vi vdd vdd d_mos L=0.18u W=0.69u
M2 1 vi 0 0 e_mos L=0.18u W=0.27u

.model d_mos pmos (KP=75u Vto=-0.5 lambda=0.02 Tox=100n, Cgso=2.288n, Cgdo=138.5p, Cbd=899.2p)
.model e_mos nmos (KP=300u Vto=0.5 lambda=0.02 Tox=100n, Cgso=73.61p, Cgdo=6.487p, Cbd=74.46p)


*analysis requests
.tran 0.1u 40u 0u 0.001u
*.TRAN 0.01ms 40ms 0ms 0.01ms
*.dc vi 0 2 0.01
.op
.probe
.end

