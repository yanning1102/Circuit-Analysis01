*circuit description
vdd vdd 0 dc 5
*vi vi 0 sin(0V 10V 60HZ)
vi vi 0 dc 2.35918
*diode model descriotion

M1 1 vi vdd vdd d_mos L=1.8u W=8.1u
M2 1 vi 0 0 e_mos L=1.8u W=2.7u

.model e_mos nmos (KP=300u Vto=0.5 lambda=0.02)
.model d_mos pmos (KP=75u Vto=-0.5 lambda=0.02)

*analysis requests
*.TRAN 0.01ms 40ms 0ms 0.01ms
.dc vi 0 5 0.01
.op
.probe
.end