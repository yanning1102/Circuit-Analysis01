
vi 1 0 dc 0
vbn 3 0 dc -5v
vgn 2 0 dc 5v
m1 1 2 0 3 aaa l=10u w=50u
.model aaa nmos(kp=20u vto=1v lambda=0)

vbp 4 0 dc 5v
vgp 5 0 dc -5v
m2 1 5 0 4 ccc l=10u w=50u
.model ccc pmos(kp=20u vto=-1v lambda=0)
.dc vi -5 5 10.001m
.probe
.end
